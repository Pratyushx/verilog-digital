module bufif1_gates(a,b,y);

input a;
input b;
output y;


bufif1 f7(y,a,b);





endmodule