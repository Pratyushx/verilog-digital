module and_gate(a,b,y);
input a;
input b;
output y;

and a1(y,a,b);

endmodule