module nor_gate(a,b,y);
input a;
input b;
output y;


nor a3(y,a,b);

endmodule