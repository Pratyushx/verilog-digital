module param_test;

parameter M=8;
parameter N=10;

initial

$display("In %m M=%0d, N=%0d",M,N);

endmodule
