module basic_gates(a,b,y);
input a;
input b;
output y;


buf a6(y,a,b);





endmodule