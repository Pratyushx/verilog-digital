module or_gate(a,b,y);
input a;
input b;
output y;

or a2(y,a,b);

endmodule