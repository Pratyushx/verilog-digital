module buf_gate(a,y);
input a;
output y;


buf a6(y,a);





endmodule