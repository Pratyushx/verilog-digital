module xor_gate(a,b,y);
input a;
input b;
output y;


xor a5(y,a,b);





endmodule