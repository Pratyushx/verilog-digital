module nand_gate(a,b,y);
input a;
input b;
output y;


nand a4(y,a,b);





endmodule